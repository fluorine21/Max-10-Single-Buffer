//Pixel writer
//Writes incomming pixels to memory
//Also packaged two pixels into one and writes them
//Should write to half of the current addr (shifted over by 1)

module pixel_writer
#(
parameter VSYNC_ACTIVE = 0
)
(
	input wire clk,
	input wire reset,//Active low, connected to system reset
	
	input wire [16:0] pixel_addr,//Incoming pixel write address
	input wire [7:0] pixel_data,//Incoming pixel data
	input wire pixel_WE,//Pixel latch
	input wire sram_ready,
	input wire pixel_vsync,
	
	output reg [15:0] sram_addr,
	output reg [15:0] sram_data,
	output sram_rw,
	output reg sram_start,//
	output reg frame_end,//Pulses when time has come to switch to sending process
	output reg error,//Signals when something has gone wrong (we see VSYNC before FFD9)
	output reg pixel_capture_reset,//Needed to reser the pixel capture module
	output reg [15:0] stop_addr//Last address written to
);



localparam PIXEL_ACTIVE = 1'b0;

reg [2:0] state;
reg [1:0] global_state;

//Holding the last data we wrote to check for a frame end
reg [15:0] sram_data_prev;


//Defining internal states
localparam [2:0] state_wait_first = 3'b000,//wait for first pixel
					  state_wait_first_end = 3'b001,//Wait for first pixel to end (WE goes low)
					  state_wait_second = 3'b010, //Wait for first pixel
					  state_end_write = 3'b011; //Wait for WE to go low, also check addr
					  
//Defining global states
localparam [1:0] state_wait_frame_end = 2'b00,//Waiting for VSYNC to go active
					  state_wait_frame = 2'b01,//Waitinf for VSYNC to turn off
					  state_frame_capture = 2'b10;//Capturing the frame
	
//Initial start_up values	
initial begin
	reset_regs();
end					  


always @ (negedge clk or negedge reset) begin
	
	if(reset == 1'b0) begin
		reset_regs();
	end
	else begin
		case (global_state)
		
			//Reset state needed to catch the frame
			state_wait_frame_end: begin
				//Reset the pixel counter.
				pixel_capture_reset <= 1'b0;
				if(pixel_vsync == VSYNC_ACTIVE)begin
					global_state <= state_wait_frame;
				end
			end
		
			//Waiting for the frame to begin
			state_wait_frame: begin
				//Reset the pixel counter.
				pixel_capture_reset <= 1'b0;
			//If the frame is starting
					if(pixel_vsync != VSYNC_ACTIVE)begin
						//Turn on pixel capture
						pixel_capture_reset <= 1'b1;
						
						//Capture the frame
						global_state <= state_frame_capture;
						//state <= state_wait_first;
						
						//Turn off our vsync
						frame_end <= 1'b0;
					end
			
			end
			
			//Writing the frame to memory
			state_frame_capture: begin
			
		
				//State machine
				case(state)
				
					state_wait_first: begin
						//If we see VSYNC active for some reason, then something has gone wrong
						if(pixel_vsync == VSYNC_ACTIVE) begin
							//Wait for the frame to start again
							global_state <= state_wait_frame;
							//Set the error flag
							error <= 1'b1;
						end
						//If we see an incomming pixel
						else if(pixel_WE == 1'b1) begin
							//Store it in the lower portion of the sram data buffer
							sram_data[7:0] <= pixel_data; 
							//store the address divided by 2 in our address buffer
							sram_addr <= (pixel_addr[15:0] >> 1);
							
							//Advance to the next state
							state <= state_wait_first_end;
						end
					
					end
					
					state_wait_first_end: begin
						//If the write has ended
						if(pixel_WE == 1'b0)begin
							//Advance to the next state
							state <= state_wait_second;
						end
					
					end
					
					state_wait_second: begin
						//If we see the second pixel
						if(pixel_WE == 1'b1) begin
							//Write the pixel to the upper half of the data buffer
							sram_data[15:8] = pixel_data;
							//If we can write to memory
							if(sram_ready == 1'b1) begin
								//Start the write process
								sram_start <= 1'b0;
							
								//Wait for the write to end
								state <= state_end_write;
							end
					
						end
					end
					
					
					state_end_write: begin
						//if pixel write went low
						sram_start <= 1'b1;
						if(pixel_WE == 1'b0) begin 
							//If the frame is done
							if(sram_data == 16'hD9FF || (sram_data[7:0] == 8'hD9 && sram_data_prev[15:8] == 8'hFF)) begin
								//Store the stop address
								stop_addr <= sram_addr;
								//Indicate that the frame has ended
								frame_end <= 1'b1;
								
								//HALT HERE until reset
								//global_state <= state_wait_frame;
								//state <= state_wait_first;
							end
							else begin
							//Store the last word
							sram_data_prev <= sram_data;
							//Reset
							state <= state_wait_first;
							end
						end		
					end
		
		
				endcase//local case
			
			end//local clause
		endcase//global case
		
	end//not reset

end//always


//Task for resetting everything
task reset_regs;
begin
	sram_addr <= 16'b0;
	sram_data <= 16'b0;
	sram_start <= 1'b1;//active low
	
	frame_end <= 1'b0;
	
	//Initializing our state
	state <= state_wait_first;
	global_state <= state_wait_frame_end;
	
	error <= 1'b0;
	
	pixel_capture_reset <= 1'b0;//Keep pixel capture in reset if we are reset
	
	//Reset the previous data register
	sram_data_prev <= 16'b0;
	
	
	stop_addr <= 16'b0;
end
endtask


assign sram_rw = 1'b0; //0 for a write

endmodule
